module PC(entrada_instrucao, saida_instrucao);
	input [31:0]entrada_instrucao;
	output [31:0]saida_instrucao;
	assign saida_instrucao = entrada_instrucao;
endmodule 