module instruction_memory(read_adress);
	input [31:0] read_adress;
	wire [4:0]read_register1, read_register2, entrada_mux2;
	wire [15:0] parte_final_da_instrucao;
endmodule 